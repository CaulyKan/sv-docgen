
module test(input wire[9:0] a [0:4], b, inout c);

endmodule

module test2(a,b,c);
    input a,c;
    wire a;
    input logic[7:0] b [3:0];
endmodule